


`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    15:11:29 11/26/2016 
// Design Name: 
// Module Name:    VRAM 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module redRAM(
	input CLK,
	input SSR,//reset here
	input EN,
	input WE,
	input [13:0] ADDR,
	input DI,
	output DO
);


		
/*
 - 16Kx1 VRAM memory(single-port) 

 - I create 3 instances of that module, one for each color
 to make the 128x96MEM
*/ 

   RAMB16_S1 #(
      .INIT(1'b0),  // Value of output RAM registers at startup
      .SRVAL(1'b0), // Output value upon SSR assertion
      .WRITE_MODE("WRITE_FIRST"), // WRITE_FIRST, READ_FIRST or NO_CHANGE

      // The following INIT_xx declarations specify the initial contents of the RAM
      // Address 0 to 4095
		/*
*************************   1st shape   ****************************************
      */		       
      .INIT_00(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),//kokkino
      .INIT_01(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),//aspro
      .INIT_02(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),//kokkino
      .INIT_03(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),//aspro
      .INIT_04(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),//...
      .INIT_05(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_06(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_07(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_08(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_09(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_0A(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
		.INIT_0B(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      /*
*************************   2nd shape   ****************************************
      */		
      .INIT_0C(256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_0D(256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_0E(256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),//...
      .INIT_0F(256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),//aspro
                         // Address 4096 to 8191
      .INIT_10(256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),//prasino
      .INIT_11(256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),//aspro
      .INIT_12(256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),//prasino
      .INIT_13(256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),//aspro
      .INIT_14(256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),//...
      .INIT_15(256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_16(256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_17(256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      /*
*************************   3rd shape   *****************************************************		
		*/
		.INIT_18(256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_19(256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_1A(256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_1B(256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_1C(256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_1D(256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_1E(256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_1F(256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),//ASPRO
      // Address 8192 to 12287
      .INIT_20(256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),//mple
      .INIT_21(256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),//aspro
      .INIT_22(256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_23(256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      /*
*************************   4th shape   ****************************************************
      (prasino-mple-aspro-aspro-aspro-kokkino)*
		        0           F           F
		*/	                                   
		.INIT_24(256'h00000000000000000000000000000000_0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0F),
      .INIT_25(256'h0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0F_0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0F),
      .INIT_26(256'h0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0F_0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0F),
      .INIT_27(256'h0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0F_0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0F),
      .INIT_28(256'h0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0F_0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0F),
      .INIT_29(256'h0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0F_0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0F),
      .INIT_2A(256'h0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0F_0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0F),
      .INIT_2B(256'h0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0F_0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0F),
      .INIT_2C(256'h0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0F_0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0F),
      .INIT_2D(256'h0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0F_0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0F),
      .INIT_2E(256'h0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0F_0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0F),
      .INIT_2F(256'h0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0F_0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0F),
      // Address 12288 to 16383
      /*
************************  END OF MEMORY  ************************************
		(prasino-mple-aspro-aspro-aspro-kokkino)*
		 00FFFF00FFFF....0000_0000_1111_1111_1111_1111_0000_0000---0_FF
		*/
		                                               
      .INIT_30(256'h000000000000000000000000000000000FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0F),//mia mavri grammi edw
      .INIT_31(256'hFF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0F),
      .INIT_32(256'hFF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0F),
      .INIT_33(256'hFF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0F),
      .INIT_34(256'hFF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0F),
      .INIT_35(256'hFF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0F),
      .INIT_36(256'hFF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0F),
      .INIT_37(256'hFF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0F),
      .INIT_38(256'hFF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0F),
      .INIT_39(256'hFF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0F),
      .INIT_3A(256'hFF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0F),
      .INIT_3B(256'hFF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0F),
      .INIT_3C(256'hFF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0F),
      .INIT_3D(256'hFF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0F),
      .INIT_3E(256'hFF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0F),
      .INIT_3F(256'hFF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0F)
   ) RAMB16 (
      .DO(DO),      // 1-bit Data Output
      .ADDR(ADDR),  // 14-bit Address Input
      .CLK(CLK),    // Clock
      .DI(DI),      // 1-bit Data Input
      .EN(EN),      // RAM Enable Input
      .SSR(SSR),    // Synchronous Set/Reset Input
      .WE(WE)       // Write Enable Input   );
   );


endmodule
